/* Copyright (C) 2017 Daniel Page <csdsp@bristol.ac.uk>
 *
 * Use of this source code is restricted per the CC BY-NC-ND license, a copy of 
 * which can be found via http://creativecommons.org (and should be included as 
 * LICENSE.txt within the associated archive or repository).
 */

module example( output wire co,
                output wire  s,

                input  wire  x,
                input  wire  y );

  xor t0(  s, x, y );
  and t1( co, x, y );

endmodule
