/* Copyright (C) 2017 Daniel Page <csdsp@bristol.ac.uk>
 *
 * Use of this source code is restricted per the CC BY-NC-ND license, a copy of 
 * which can be found via http://creativecommons.org (and should be included as 
 * LICENSE.txt within the associated archive or repository).
 */

module add_4bit( output wire           co,
                 output wire [ 3 : 0 ] r,

                  input wire           ci,
                  input wire [ 3 : 0 ] x,
                  input wire [ 3 : 0 ] y );

endmodule
