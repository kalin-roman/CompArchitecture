/* Copyright (C) 2017 Daniel Page <csdsp@bristol.ac.uk>
 *
 * Use of this source code is restricted per the CC BY-NC-ND license, a copy of 
 * which can be found via http://creativecommons.org (and should be included as 
 * LICENSE.txt within the associated archive or repository).
 */

module ctr_4bit_fflop(  input wire           mode,
                        input wire           rst,

                        input wire           clk,

                       output wire [ 3 : 0 ] r );

endmodule
